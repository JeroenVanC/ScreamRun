module score_counter (display_col, display_row, reset, visible, clock, hit, score_red, score_green, score_blue, score_visible);
